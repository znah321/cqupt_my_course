library verilog;
use verilog.vl_types.all;
entity dMogan_Bool_2_vlg_vec_tst is
end dMogan_Bool_2_vlg_vec_tst;
