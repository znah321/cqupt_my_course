library verilog;
use verilog.vl_types.all;
entity MUX151_vlg_vec_tst is
end MUX151_vlg_vec_tst;
