library verilog;
use verilog.vl_types.all;
entity Scan_Module_vlg_vec_tst is
end Scan_Module_vlg_vec_tst;
