library verilog;
use verilog.vl_types.all;
entity RS_Latch_vlg_check_tst is
    port(
        Reset           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end RS_Latch_vlg_check_tst;
