library verilog;
use verilog.vl_types.all;
entity Buzzer_Hour_Simulation_vlg_vec_tst is
end Buzzer_Hour_Simulation_vlg_vec_tst;
