library verilog;
use verilog.vl_types.all;
entity Second_Count_vlg_vec_tst is
end Second_Count_vlg_vec_tst;
