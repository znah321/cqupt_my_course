library verilog;
use verilog.vl_types.all;
entity four_xorGate_vlg_vec_tst is
end four_xorGate_vlg_vec_tst;
