library verilog;
use verilog.vl_types.all;
entity block1_vlg_vec_tst is
end block1_vlg_vec_tst;
