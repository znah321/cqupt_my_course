library verilog;
use verilog.vl_types.all;
entity andGate_vlg_vec_tst is
end andGate_vlg_vec_tst;
