library verilog;
use verilog.vl_types.all;
entity xxx is
    port(
        pin_name2       : out    vl_logic;
        pin_name1       : in     vl_logic
    );
end xxx;
