library verilog;
use verilog.vl_types.all;
entity TimingModule_Second_Minute_vlg_sample_tst is
    port(
        Input           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end TimingModule_Second_Minute_vlg_sample_tst;
