library verilog;
use verilog.vl_types.all;
entity Buzzer_Clock_Simulation_vlg_check_tst is
    port(
        Buzzer          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Buzzer_Clock_Simulation_vlg_check_tst;
