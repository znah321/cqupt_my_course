library verilog;
use verilog.vl_types.all;
entity RS_Latch_vlg_vec_tst is
end RS_Latch_vlg_vec_tst;
