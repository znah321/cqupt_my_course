library verilog;
use verilog.vl_types.all;
entity counter_vlg_vec_tst is
end counter_vlg_vec_tst;
