library verilog;
use verilog.vl_types.all;
entity Timing_Module_vlg_sample_tst is
    port(
        Input           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Timing_Module_vlg_sample_tst;
