library verilog;
use verilog.vl_types.all;
entity block2_vlg_check_tst is
    port(
        G               : in     vl_logic;
        R               : in     vl_logic;
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end block2_vlg_check_tst;
