library verilog;
use verilog.vl_types.all;
entity Count_Second_vlg_vec_tst is
end Count_Second_vlg_vec_tst;
