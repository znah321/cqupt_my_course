library verilog;
use verilog.vl_types.all;
entity notGate_vlg_vec_tst is
end notGate_vlg_vec_tst;
