library verilog;
use verilog.vl_types.all;
entity Count_Hour_vlg_vec_tst is
end Count_Hour_vlg_vec_tst;
