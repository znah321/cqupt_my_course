library verilog;
use verilog.vl_types.all;
entity D_trigger_vlg_vec_tst is
end D_trigger_vlg_vec_tst;
