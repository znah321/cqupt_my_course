library verilog;
use verilog.vl_types.all;
entity Test_vlg_vec_tst is
end Test_vlg_vec_tst;
