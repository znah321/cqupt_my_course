library verilog;
use verilog.vl_types.all;
entity Timing_Module_vlg_vec_tst is
end Timing_Module_vlg_vec_tst;
