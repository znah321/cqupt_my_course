library verilog;
use verilog.vl_types.all;
entity xorGate_vlg_vec_tst is
end xorGate_vlg_vec_tst;
