library verilog;
use verilog.vl_types.all;
entity Count_S_vlg_vec_tst is
end Count_S_vlg_vec_tst;
