library verilog;
use verilog.vl_types.all;
entity Bit_Selective_Signal_Generator_vlg_sample_tst is
    port(
        Clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Bit_Selective_Signal_Generator_vlg_sample_tst;
