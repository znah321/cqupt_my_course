library verilog;
use verilog.vl_types.all;
entity notGate_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end notGate_vlg_sample_tst;
