library verilog;
use verilog.vl_types.all;
entity dMogan_Bool_1_vlg_check_tst is
    port(
        YLeft           : in     vl_logic;
        YRight          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end dMogan_Bool_1_vlg_check_tst;
