library verilog;
use verilog.vl_types.all;
entity xnorGate_logicgate_vlg_vec_tst is
end xnorGate_logicgate_vlg_vec_tst;
