library verilog;
use verilog.vl_types.all;
entity Count_Hour_vlg_sample_tst is
    port(
        Clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Count_Hour_vlg_sample_tst;
