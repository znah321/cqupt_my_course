library verilog;
use verilog.vl_types.all;
entity mux3_en_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux3_en_vlg_check_tst;
