library verilog;
use verilog.vl_types.all;
entity block2_vlg_check_tst is
    port(
        EB              : in     vl_logic;
        GB              : in     vl_logic;
        LB              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end block2_vlg_check_tst;
