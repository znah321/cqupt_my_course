library verilog;
use verilog.vl_types.all;
entity compare_gate_vlg_vec_tst is
end compare_gate_vlg_vec_tst;
