library verilog;
use verilog.vl_types.all;
entity lab3_vlg_sample_tst is
    port(
        CP              : in     vl_logic;
        en              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab3_vlg_sample_tst;
