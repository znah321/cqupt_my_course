library verilog;
use verilog.vl_types.all;
entity TimingModule_Second_Minute_vlg_vec_tst is
end TimingModule_Second_Minute_vlg_vec_tst;
