library verilog;
use verilog.vl_types.all;
entity Buzzer_Clock_Simulation_vlg_vec_tst is
end Buzzer_Clock_Simulation_vlg_vec_tst;
