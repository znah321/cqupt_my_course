library verilog;
use verilog.vl_types.all;
entity mux3_vlg_vec_tst is
end mux3_vlg_vec_tst;
