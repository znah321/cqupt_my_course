library verilog;
use verilog.vl_types.all;
entity mux3_en_vlg_vec_tst is
end mux3_en_vlg_vec_tst;
