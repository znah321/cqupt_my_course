library verilog;
use verilog.vl_types.all;
entity Buzzer_Hour_Simulation_vlg_check_tst is
    port(
        Buzzer          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Buzzer_Hour_Simulation_vlg_check_tst;
