library verilog;
use verilog.vl_types.all;
entity or_not_Gate_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end or_not_Gate_vlg_check_tst;
