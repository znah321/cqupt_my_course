library verilog;
use verilog.vl_types.all;
entity dMogan_Bool_2_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end dMogan_Bool_2_vlg_check_tst;
