library verilog;
use verilog.vl_types.all;
entity xxx_vlg_vec_tst is
end xxx_vlg_vec_tst;
