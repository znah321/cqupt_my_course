library verilog;
use verilog.vl_types.all;
entity orGate_vlg_vec_tst is
end orGate_vlg_vec_tst;
