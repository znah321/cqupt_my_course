library verilog;
use verilog.vl_types.all;
entity DigitalClock_vlg_vec_tst is
end DigitalClock_vlg_vec_tst;
