library verilog;
use verilog.vl_types.all;
entity or_not_Gate_vlg_vec_tst is
end or_not_Gate_vlg_vec_tst;
