library verilog;
use verilog.vl_types.all;
entity block2_vlg_vec_tst is
end block2_vlg_vec_tst;
