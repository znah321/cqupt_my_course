library verilog;
use verilog.vl_types.all;
entity lab4_vlg_sample_tst is
    port(
        CP              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab4_vlg_sample_tst;
