library verilog;
use verilog.vl_types.all;
entity four_andGate_vlg_vec_tst is
end four_andGate_vlg_vec_tst;
