library verilog;
use verilog.vl_types.all;
entity TimeingModule_Minute_Hour_vlg_vec_tst is
end TimeingModule_Minute_Hour_vlg_vec_tst;
